library verilog;
use verilog.vl_types.all;
entity pipeCPU_vlg_tst is
end pipeCPU_vlg_tst;
